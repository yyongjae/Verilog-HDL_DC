module ex01(in1,in2,out1);
    input in1, in2;
    output out1;
    wire in1, in2;
    wire out1;
    assign out1 = in1 & in2;
endmodule